library IEEE;
use IEEE.std_logic_1164.all;

package bus_6digit is
	type bus_array is array(0 to 5) of std_logic_vector(5 downto 0);
end package bus_6digit;